../clk/rt_clk.vhdl