-- file : lfsr4.vhdl
-- parameterised LFSR generator
-- data from http://www.physics.otago.ac.nz/px/research/electronics/papers/technical-reports/lfsr_table.pdf
-- version oct. 8 01:09:20 CEST 2010
-- Copyright (C) 2010 Yann GUIDON
--
-- This program is free software: you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation, either version 3 of the License, or
-- (at your option) any later version.
--
-- This program is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
--
-- You should have received a copy of the GNU General Public License
-- along with this program.  If not, see <http://www.gnu.org/licenses/>.

library ieee;
use ieee.std_logic_1164.all;

entity lfsr4 is
  generic(
    size : integer := 8
  );
  port(
    clk, reset, din : in std_logic := '0';
    lfsr : inout std_ulogic_vector(size downto 1);
    init_val : in std_ulogic_vector(size downto 1) := (1=>'1', others=>'0'); -- leave "open" or connect to a constant only
    s : out std_logic
  );
end lfsr4;

architecture fibonacci of lfsr4 is
  constant first_poly : integer := 5;
  constant  last_poly : integer := 786;

  type poly_array_type is array(first_poly to last_poly, 0 to 2) of integer;
  constant poly4_array : poly_array_type := (
(4, 3, 2),
(5, 3, 2),
(6, 5, 4),
(6, 5, 4),
(8, 6, 5),
(9, 7, 6),
(10, 9, 7),
(11, 8, 6),
(12, 10, 9),
(13, 11, 9),
(14, 13, 11),
(14, 13, 11),
(16, 15, 14),
(17, 16, 13),
(18, 17, 14),
(19, 16, 14),
(20, 19, 16),
(19, 18, 17),
(22, 20, 18),
(23, 21, 20),
(24, 23, 22),
(25, 24, 20),
(26, 25, 22),
(27, 24, 22),
(28, 27, 25),
(29, 26, 24),
(30, 29, 28),
(30, 26, 25),
(32, 29, 27),
(31, 30, 26),
(34, 28, 27),
(35, 29, 28),
(36, 33, 31),
(37, 33, 32),
(38, 35, 32),
(37, 36, 35),
(40, 39, 38),
(40, 37, 35),
(42, 38, 37),
(42, 39, 38),
(44, 42, 41),
(40, 39, 38),
(46, 43, 42),
(44, 41, 39),
(45, 44, 43),
(48, 47, 46),
(50, 48, 45),
(51, 49, 46),
(52, 51, 47),
(51, 48, 46),
(54, 53, 49),
(54, 52, 49),
(55, 54, 52),
(57, 53, 52),
(57, 55, 52),
(58, 56, 55),
(60, 59, 56),
(59, 57, 56),
(62, 59, 58),
(63, 61, 60),
(64, 62, 61),
(60, 58, 57),
(66, 65, 62),
(67, 63, 61),
(67, 64, 63),
(69, 67, 65),
(70, 68, 66),
(69, 63, 62),
(71, 70, 69),
(71, 70, 67),
(74, 72, 69),
(74, 72, 71),
(75, 72, 71),
(77, 76, 71),
(77, 76, 75),
(78, 76, 71),
(79, 78, 75),
(78, 76, 73),
(81, 79, 76),
(83, 77, 75),
(84, 83, 77),
(84, 81, 80),
(86, 82, 80),
(80, 79, 77),
(86, 84, 83),
(88, 87, 85),
(90, 86, 83),
(90, 87, 86),
(91, 90, 87),
(93, 89, 88),
(94, 90, 88),
(90, 87, 86),
(95, 93, 91),
(97, 91, 90),
(95, 94, 92),
(98, 93, 92),
(100, 95, 94),
(99, 97, 96),
(102, 99, 94),
(103, 94, 93),
(104, 99, 98),
(105, 101, 100),
(105, 99, 98),
(103, 97, 96),
(107, 105, 104),
(109, 106, 104),
(109, 107, 104),
(108, 106, 101),
(111, 110, 108),
(113, 112, 103),
(110, 108, 107),
(114, 111, 110),
(116, 115, 112),
(116, 113, 112),
(116, 111, 110),
(118, 114, 111),
(120, 116, 113),
(121, 120, 116),
(122, 119, 115),
(119, 118, 117),
(120, 119, 118),
(124, 122, 119),
(126, 124, 120),
(127, 126, 121),
(128, 125, 124),
(129, 128, 125),
(129, 128, 123),
(130, 127, 123),
(131, 125, 124),
(133, 129, 127),
(132, 131, 129),
(134, 133, 128),
(136, 133, 126),
(137, 131, 130),
(136, 134, 131),
(139, 136, 132),
(140, 135, 128),
(141, 139, 132),
(141, 140, 138),
(142, 140, 137),
(144, 140, 139),
(144, 143, 141),
(145, 143, 136),
(145, 143, 141),
(142, 140, 139),
(148, 147, 142),
(150, 149, 148),
(150, 149, 146),
(149, 148, 145),
(153, 149, 145),
(151, 150, 148),
(153, 151, 147),
(155, 152, 151),
(153, 152, 150),
(156, 153, 148),
(158, 157, 155),
(159, 158, 155),
(158, 155, 154),
(160, 157, 156),
(159, 158, 152),
(162, 157, 156),
(164, 163, 156),
(165, 163, 161),
(162, 159, 152),
(164, 163, 161),
(169, 166, 161),
(169, 166, 165),
(169, 165, 161),
(171, 168, 165),
(169, 166, 165),
(173, 171, 169),
(167, 165, 164),
(175, 174, 172),
(176, 171, 170),
(178, 177, 175),
(173, 170, 168),
(180, 175, 174),
(181, 176, 174),
(179, 176, 175),
(177, 176, 175),
(184, 182, 177),
(180, 178, 177),
(182, 181, 180),
(186, 183, 182),
(187, 184, 183),
(188, 184, 177),
(187, 185, 184),
(190, 178, 177),
(189, 186, 184),
(192, 191, 190),
(193, 192, 187),
(194, 187, 185),
(195, 193, 188),
(193, 190, 183),
(198, 195, 190),
(198, 197, 195),
(199, 198, 195),
(198, 196, 195),
(202, 196, 195),
(201, 200, 194),
(203, 200, 196),
(201, 197, 196),
(206, 201, 198),
(207, 205, 199),
(207, 206, 204),
(207, 206, 198),
(203, 201, 200),
(209, 208, 205),
(211, 208, 207),
(213, 211, 209),
(212, 210, 209),
(215, 213, 209),
(213, 212, 211),
(217, 211, 210),
(218, 215, 211),
(211, 210, 208),
(219, 215, 213),
(220, 217, 214),
(221, 219, 218),
(222, 217, 212),
(224, 220, 215),
(223, 219, 216),
(223, 218, 217),
(226, 217, 216),
(228, 225, 219),
(224, 223, 222),
(229, 227, 224),
(228, 223, 221),
(232, 229, 224),
(232, 225, 223),
(234, 229, 226),
(229, 228, 226),
(236, 233, 230),
(237, 236, 233),
(238, 232, 227),
(237, 235, 232),
(237, 233, 232),
(241, 236, 231),
(242, 238, 235),
(243, 240, 235),
(244, 241, 239),
(245, 244, 235),
(245, 243, 238),
(238, 234, 233),
(248, 245, 242),
(247, 245, 240),
(249, 247, 244),
(251, 247, 241),
(252, 247, 246),
(253, 252, 247),
(253, 252, 250),
(254, 251, 246),
(255, 251, 250),
(254, 252, 249),
(257, 253, 249),
(253, 252, 250),
(257, 255, 254),
(258, 254, 253),
(261, 258, 252),
(263, 255, 254),
(263, 262, 260),
(265, 260, 259),
(264, 261, 259),
(267, 264, 258),
(268, 263, 262),
(267, 263, 260),
(265, 264, 260),
(270, 266, 263),
(272, 271, 266),
(272, 267, 265),
(266, 265, 264),
(275, 273, 270),
(274, 271, 265),
(277, 274, 273),
(278, 275, 274),
(278, 275, 271),
(280, 277, 272),
(278, 277, 272),
(278, 276, 271),
(279, 278, 276),
(280, 278, 275),
(285, 276, 271),
(285, 282, 281),
(287, 278, 277),
(286, 285, 277),
(288, 287, 285),
(286, 280, 279),
(291, 289, 285),
(292, 287, 282),
(292, 291, 285),
(293, 291, 290),
(292, 287, 285),
(296, 293, 292),
(294, 290, 287),
(295, 293, 288),
(290, 288, 287),
(299, 296, 292),
(297, 293, 290),
(297, 291, 290),
(303, 302, 293),
(303, 299, 298),
(305, 303, 299),
(305, 303, 299),
(306, 299, 293),
(307, 302, 299),
(309, 305, 302),
(308, 306, 304),
(307, 302, 301),
(312, 310, 306),
(311, 305, 300),
(314, 306, 305),
(309, 305, 304),
(315, 313, 310),
(313, 312, 310),
(318, 317, 308),
(319, 317, 316),
(319, 316, 314),
(321, 320, 305),
(322, 320, 313),
(321, 320, 318),
(323, 320, 315),
(325, 323, 316),
(325, 322, 319),
(323, 321, 319),
(326, 323, 321),
(328, 323, 322),
(329, 325, 321),
(325, 321, 320),
(331, 329, 325),
(333, 330, 327),
(333, 328, 325),
(335, 332, 329),
(336, 331, 327),
(336, 335, 332),
(332, 329, 323),
(337, 336, 329),
(336, 330, 327),
(341, 340, 331),
(338, 335, 333),
(338, 334, 333),
(343, 341, 337),
(344, 339, 335),
(344, 337, 336),
(344, 341, 340),
(347, 344, 343),
(340, 337, 336),
(348, 345, 343),
(346, 341, 339),
(349, 346, 344),
(349, 341, 340),
(354, 350, 349),
(349, 347, 346),
(355, 347, 346),
(351, 350, 344),
(358, 352, 350),
(359, 335, 334),
(360, 357, 354),
(360, 351, 344),
(362, 356, 355),
(363, 359, 352),
(360, 359, 356),
(362, 359, 352),
(365, 363, 358),
(361, 359, 351),
(367, 359, 358),
(368, 367, 365),
(369, 368, 363),
(369, 365, 357),
(371, 366, 365),
(369, 368, 366),
(374, 368, 367),
(371, 369, 368),
(376, 374, 369),
(374, 365, 363),
(375, 370, 369),
(377, 374, 366),
(380, 379, 376),
(379, 375, 364),
(382, 378, 374),
(378, 369, 368),
(383, 381, 379),
(381, 380, 376),
(385, 379, 378),
(387, 385, 374),
(384, 380, 379),
(388, 380, 377),
(390, 389, 385),
(386, 382, 379),
(392, 391, 386),
(392, 387, 386),
(390, 389, 384),
(392, 390, 389),
(392, 387, 385),
(393, 392, 384),
(397, 390, 388),
(398, 397, 395),
(399, 392, 389),
(399, 398, 393),
(398, 395, 394),
(400, 398, 397),
(398, 397, 388),
(402, 397, 393),
(402, 400, 398),
(407, 403, 401),
(406, 404, 402),
(407, 406, 400),
(408, 401, 399),
(409, 404, 401),
(407, 406, 403),
(405, 401, 398),
(413, 411, 406),
(414, 411, 407),
(416, 414, 407),
(417, 415, 403),
(415, 414, 404),
(412, 410, 407),
(419, 417, 416),
(421, 416, 412),
(420, 418, 414),
(422, 417, 415),
(422, 421, 418),
(415, 414, 412),
(422, 421, 416),
(426, 425, 417),
(422, 421, 419),
(419, 417, 415),
(430, 428, 426),
(429, 428, 419),
(430, 428, 422),
(429, 423, 422),
(430, 426, 423),
(432, 431, 430),
(436, 435, 431),
(436, 432, 421),
(437, 436, 431),
(439, 437, 436),
(440, 433, 430),
(440, 437, 435),
(442, 437, 433),
(435, 432, 431),
(441, 439, 438),
(442, 439, 431),
(446, 441, 438),
(444, 442, 437),
(446, 440, 438),
(443, 438, 434),
(450, 441, 435),
(448, 447, 446),
(449, 447, 438),
(449, 445, 444),
(453, 449, 444),
(454, 445, 433),
(454, 449, 446),
(453, 448, 445),
(457, 454, 447),
(459, 455, 451),
(460, 455, 454),
(457, 451, 450),
(456, 455, 452),
(460, 455, 441),
(463, 462, 457),
(460, 455, 452),
(466, 461, 456),
(464, 459, 453),
(467, 464, 460),
(468, 462, 461),
(469, 468, 465),
(470, 469, 461),
(470, 467, 465),
(465, 463, 456),
(471, 467, 466),
(475, 468, 466),
(470, 462, 461),
(477, 474, 472),
(475, 472, 470),
(473, 467, 464),
(480, 472, 471),
(477, 476, 473),
(479, 477, 474),
(483, 482, 470),
(479, 469, 468),
(481, 478, 472),
(485, 483, 478),
(487, 485, 484),
(484, 483, 480),
(485, 483, 481),
(488, 485, 480),
(491, 485, 484),
(490, 488, 483),
(493, 489, 481),
(494, 486, 480),
(494, 491, 480),
(493, 488, 486),
(495, 489, 487),
(494, 493, 488),
(499, 494, 490),
(499, 497, 496),
(498, 497, 494),
(502, 501, 500),
(502, 490, 483),
(500, 497, 493),
(501, 494, 491),
(504, 501, 494),
(505, 500, 495),
(506, 502, 501),
(501, 500, 498),
(509, 503, 501),
(510, 507, 504),
(505, 503, 500),
(511, 509, 507),
(511, 508, 501),
(514, 511, 509),
(515, 507, 505),
(516, 515, 507),
(517, 511, 507),
(509, 507, 503),
(519, 514, 512),
(518, 509, 507),
(521, 517, 510),
(523, 519, 515),
(524, 521, 519),
(525, 521, 517),
(526, 520, 518),
(526, 522, 517),
(528, 525, 522),
(527, 523, 520),
(529, 525, 519),
(529, 528, 522),
(531, 530, 529),
(533, 529, 527),
(533, 529, 527),
(533, 531, 529),
(536, 535, 527),
(537, 536, 533),
(535, 534, 529),
(537, 534, 529),
(537, 531, 528),
(540, 539, 533),
(538, 536, 532),
(538, 535, 531),
(539, 537, 532),
(545, 544, 538),
(543, 540, 534),
(545, 543, 538),
(546, 545, 533),
(546, 533, 529),
(550, 547, 542),
(550, 547, 532),
(550, 549, 542),
(551, 546, 543),
(551, 546, 545),
(549, 546, 540),
(552, 551, 550),
(553, 549, 544),
(557, 552, 550),
(554, 551, 549),
(558, 552, 550),
(560, 558, 551),
(561, 554, 549),
(563, 561, 558),
(564, 559, 554),
(564, 561, 560),
(563, 557, 556),
(558, 557, 551),
(568, 559, 557),
(563, 558, 552),
(569, 566, 561),
(571, 564, 560),
(569, 567, 563),
(569, 565, 560),
(572, 570, 569),
(573, 572, 563),
(575, 574, 569),
(562, 556, 555),
(572, 570, 567),
(579, 576, 574),
(575, 574, 568),
(579, 576, 571),
(581, 577, 575),
(581, 571, 570),
(583, 582, 577),
(584, 581, 579),
(586, 581, 576),
(577, 572, 571),
(586, 585, 579),
(588, 587, 578),
(587, 585, 582),
(591, 573, 568),
(588, 585, 584),
(586, 584, 583),
(594, 593, 586),
(592, 591, 590),
(588, 585, 583),
(597, 592, 591),
(593, 591, 590),
(599, 590, 589),
(600, 597, 589),
(596, 594, 591),
(600, 599, 597),
(600, 598, 589),
(600, 598, 595),
(602, 599, 591),
(600, 598, 595),
(606, 602, 585),
(601, 600, 597),
(602, 600, 599),
(609, 607, 601),
(607, 602, 598),
(609, 603, 594),
(613, 612, 607),
(614, 609, 608),
(614, 602, 597),
(612, 608, 607),
(615, 604, 598),
(614, 611, 610),
(619, 618, 611),
(616, 615, 609),
(612, 610, 605),
(614, 613, 612),
(617, 615, 612),
(620, 617, 613),
(623, 621, 613),
(622, 617, 613),
(626, 617, 616),
(627, 624, 623),
(628, 626, 623),
(625, 623, 617),
(629, 619, 613),
(632, 631, 626),
(631, 629, 627),
(631, 625, 621),
(632, 628, 623),
(636, 628, 623),
(637, 633, 632),
(636, 635, 629),
(638, 637, 626),
(640, 636, 622),
(636, 633, 632),
(641, 640, 632),
(634, 633, 632),
(641, 637, 634),
(635, 634, 633),
(646, 643, 642),
(647, 626, 625),
(648, 644, 638),
(644, 635, 632),
(646, 638, 637),
(647, 643, 641),
(646, 645, 643),
(649, 643, 640),
(653, 639, 638),
(646, 638, 637),
(656, 650, 649),
(651, 648, 646),
(657, 655, 644),
(657, 656, 648),
(657, 650, 649),
(659, 656, 650),
(655, 652, 649),
(662, 660, 649),
(661, 659, 654),
(664, 659, 656),
(664, 660, 649),
(658, 656, 651),
(667, 665, 664),
(669, 665, 664),
(669, 665, 662),
(667, 666, 661),
(666, 664, 663),
(671, 665, 660),
(674, 672, 669),
(675, 671, 664),
(674, 673, 669),
(675, 673, 663),
(676, 667, 661),
(679, 650, 645),
(678, 672, 670),
(681, 679, 675),
(682, 677, 672),
(681, 671, 666),
(684, 682, 681),
(684, 674, 673),
(682, 675, 673),
(682, 674, 669),
(686, 683, 681),
(687, 683, 680),
(689, 685, 678),
(687, 686, 678),
(691, 685, 678),
(691, 681, 677),
(694, 691, 686),
(694, 686, 673),
(689, 685, 681),
(690, 689, 688),
(698, 689, 684),
(698, 695, 694),
(699, 697, 685),
(701, 699, 695),
(702, 696, 691),
(701, 699, 692),
(704, 698, 697),
(697, 695, 692),
(702, 699, 692),
(706, 704, 703),
(708, 706, 705),
(709, 696, 695),
(704, 703, 700),
(709, 708, 707),
(706, 703, 696),
(709, 707, 701),
(714, 711, 708),
(706, 705, 704),
(716, 710, 701),
(717, 716, 713),
(711, 710, 707),
(718, 712, 709),
(720, 713, 712),
(721, 718, 707),
(717, 710, 707),
(719, 716, 711),
(720, 719, 716),
(725, 722, 721),
(721, 719, 716),
(726, 725, 724),
(726, 724, 718),
(726, 715, 711),
(729, 725, 723),
(729, 728, 725),
(731, 726, 725),
(724, 721, 720),
(733, 728, 727),
(730, 728, 723),
(736, 733, 732),
(730, 729, 727),
(731, 723, 721),
(737, 728, 716),
(738, 733, 732),
(741, 738, 730),
(742, 731, 730),
(743, 733, 731),
(740, 738, 737),
(738, 733, 728),
(743, 741, 737),
(744, 743, 733),
(748, 743, 742),
(746, 741, 734),
(750, 748, 740),
(749, 732, 731),
(748, 745, 740),
(742, 740, 735),
(754, 745, 743),
(755, 747, 740),
(756, 751, 750),
(757, 746, 741),
(757, 756, 750),
(757, 747, 734),
(760, 759, 758),
(761, 755, 745),
(754, 749, 747),
(761, 759, 758),
(760, 755, 754),
(757, 747, 744),
(763, 760, 759),
(764, 751, 749),
(763, 762, 760),
(768, 765, 756),
(765, 756, 754),
(767, 766, 764),
(767, 765, 763),
(767, 760, 758),
(771, 769, 768),
(773, 764, 759),
(776, 767, 761),
(775, 762, 759),
(776, 771, 769),
(775, 772, 764),
(779, 765, 764),
(780, 779, 773),
(782, 776, 773),
(778, 775, 771),
(780, 776, 775),
(782, 780, 771));

begin
  process (clk, reset)
  begin
    if reset = '1' then
      lfsr <= init_val;
    else
      if rising_edge(clk) then
        lfsr(1) <= lfsr(size)
                  xor lfsr(poly4_array(size,0))
                  xor lfsr(poly4_array(size,1))
                  xor lfsr(poly4_array(size,2))
                  xor din;
        lfsr(size downto 2) <= lfsr(size-1 downto 1);
      end if;
    end if;
  end process;

  s <= lfsr(1);
end fibonacci;
