../fb/fb_ghdl.vhdl